/*module mem_access_test(
	input
	output
	);
	wire clk, rst;
	reg createdump, wr, rd;
	reg[15:0] addr, data_in;
	
	four_bank_mem memory0 (.clk (clk), .rst (rst), .createdump (createdump), .addr (mem_addr), .data_in (mem_in), .wr (memwr), .rd (memrd), .data_out (mem_out), .stall (mem_stall), .busy (mem_busy), .err (mem_err));
	clkrst clkgen (.clk (clk), .rst (rst), .err(1'b0));




 
endmodule */
